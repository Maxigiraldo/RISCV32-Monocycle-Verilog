module Control_Unit (
   input [6:0] opcode,
   input [2:0] funct3,
   input [6:0] funct7,
   output reg branch,
   output reg mem_read,
   output reg mem_to_reg,
   output reg [1:0] alu_op,
   output reg mem_write,
   output reg alu_src,
   output reg reg_write
);

   always @(*) begin
       // Valores por defecto
       {branch, mem_read, mem_to_reg, mem_write, alu_src, reg_write} = 6'b0;
       alu_op = 2'b00;
       
       case (opcode)
           7'b0110011: begin // R-type
               reg_write = 1;
               alu_op = 2'b10;
           end
           
           7'b0010011: begin // I-type (ALU)
               alu_src = 1;
               reg_write = 1;
               alu_op = 2'b10;
           end
           
           7'b0000011: begin // Load
               alu_src = 1;
               mem_to_reg = 1;
               reg_write = 1;
               mem_read = 1;
               alu_op = 2'b00;
           end
           
           7'b0100011: begin // Store
               alu_src = 1;
               mem_write = 1;
               alu_op = 2'b00;
           end
           
           7'b1100011: begin // Branch
               branch = 1;
               alu_op = 2'b01;
           end
			  
			  default: begin
               // NOP o instrucción no reconocida
               {branch, mem_read, mem_to_reg, mem_write, alu_src, reg_write} = 6'b0;
               alu_op = 2'b00;
           end
       endcase
   end

endmodule
